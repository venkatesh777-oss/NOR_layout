magic
tech scmos
timestamp 1764002479
<< nwell >>
rect -17 4 28 19
<< polysilicon >>
rect -6 18 -2 20
rect 10 18 14 20
rect -6 -5 -2 5
rect 10 3 14 5
rect 3 -2 14 3
rect -13 -10 -2 -5
rect -6 -18 -2 -10
rect 10 -18 14 -2
rect -6 -33 -2 -31
rect 10 -33 14 -31
<< ndiffusion >>
rect -15 -31 -6 -18
rect -2 -31 10 -18
rect 14 -31 27 -18
<< pdiffusion >>
rect -15 5 -6 18
rect -2 5 10 18
rect 14 5 27 18
<< metal1 >>
rect -16 31 26 36
rect -14 7 -7 31
rect 17 -4 24 15
rect 0 -11 37 -4
rect -14 -41 -7 -21
rect 0 -29 7 -11
rect 18 -41 25 -21
rect -15 -46 27 -41
<< ntransistor >>
rect -6 -31 -2 -18
rect 10 -31 14 -18
<< ptransistor >>
rect -6 5 -2 18
rect 10 5 14 18
<< labels >>
rlabel metal1 17 -11 37 -4 1 out
rlabel metal1 -7 31 19 35 5 vdd
rlabel metal1 -4 -46 22 -42 1 gnd
rlabel polysilicon 3 -2 14 3 1 b
rlabel polysilicon -13 -10 -2 -5 1 a
<< end >>
